`define ENABLE_XILINX_PRIMITIVES
